* C:\Users\Lucas.ordinateur\Documents\PPE\pr�sentation\schemas pspice\debitmetre potentiometre raz\schema.sch

* Schematics Version 9.1 - Web Update 1
* Sun Apr 08 11:03:54 2012



** Analysis setup **
.tran 100ns 100ms 0 10ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "schema.net"
.INC "schema.als"


.probe


.END
